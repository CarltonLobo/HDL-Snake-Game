`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/27/2025 11:32:54 AM
// Design Name: 
// Module Name: welcome_by8
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module welcome_by8
	(
		input wire clk,
		input wire [5:0] row,
		input wire [6:0] col,
		input wire [1:0] mode,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [6:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		13'b0010100001100: color_data = 12'b010010101111;
		13'b0010100010000: color_data = 12'b010010101111;
		13'b0010100010011: color_data = 12'b010010101111;
		13'b0010100010100: color_data = 12'b010010101111;
		13'b0010100010101: color_data = 12'b010010101111;
		13'b0010100010110: color_data = 12'b010010101111;
		13'b0010100011000: color_data = 12'b010010101111;
		13'b0010100011111: color_data = 12'b010010101111;
		13'b0010100100000: color_data = 12'b010010101111;
		13'b0010100100001: color_data = 12'b010010101111;
		13'b0010100100100: color_data = 12'b010010101111;
		13'b0010100100101: color_data = 12'b010010101111;
		13'b0010100100110: color_data = 12'b010010101111;
		13'b0010100101001: color_data = 12'b010010101111;
		13'b0010100101101: color_data = 12'b010010101111;
		13'b0010100110000: color_data = 12'b010010101111;
		13'b0010100110001: color_data = 12'b010010101111;
		13'b0010100110010: color_data = 12'b010010101111;
		13'b0010100110011: color_data = 12'b010010101111;
		13'b0010100111001: color_data = 12'b010010101111;
		13'b0010100111010: color_data = 12'b010010101111;
		13'b0010100111011: color_data = 12'b010010101111;
		13'b0010100111100: color_data = 12'b010010101111;
		13'b0010100111101: color_data = 12'b010010101111;
		13'b0010101000000: color_data = 12'b010010101111;
		13'b0010101000001: color_data = 12'b010010101111;
		13'b0010101000010: color_data = 12'b010010101111;

		13'b0010110001100: color_data = 12'b010010101111;
		13'b0010110010000: color_data = 12'b010010101111;
		13'b0010110010010: color_data = 12'b010010101111;
		13'b0010110010011: color_data = 12'b010010101111;
		13'b0010110011000: color_data = 12'b010010101111;
		13'b0010110011110: color_data = 12'b010010101111;
		13'b0010110011111: color_data = 12'b010010101111;
		13'b0010110100100: color_data = 12'b010010101111;
		13'b0010110100110: color_data = 12'b010010101111;
		13'b0010110101001: color_data = 12'b010010101111;
		13'b0010110101010: color_data = 12'b010010101111;
		13'b0010110101100: color_data = 12'b010010101111;
		13'b0010110101101: color_data = 12'b010010101111;
		13'b0010110101111: color_data = 12'b010010101111;
		13'b0010110110000: color_data = 12'b010010101111;
		13'b0010110111011: color_data = 12'b010010101111;
		13'b0010111000000: color_data = 12'b010010101111;
		13'b0010111000010: color_data = 12'b010010101111;

		13'b0011000001100: color_data = 12'b010010101111;
		13'b0011000010000: color_data = 12'b010010101111;
		13'b0011000010010: color_data = 12'b010010101111;
		13'b0011000010011: color_data = 12'b010010101111;
		13'b0011000011000: color_data = 12'b010010101111;
		13'b0011000011101: color_data = 12'b010010101111;
		13'b0011000011110: color_data = 12'b010010101111;
		13'b0011000100011: color_data = 12'b010010101111;
		13'b0011000100111: color_data = 12'b010010101111;
		13'b0011000101001: color_data = 12'b010010101111;
		13'b0011000101010: color_data = 12'b010010101111;
		13'b0011000101100: color_data = 12'b010010101111;
		13'b0011000101101: color_data = 12'b010010101111;
		13'b0011000101111: color_data = 12'b010010101111;
		13'b0011000110000: color_data = 12'b010010101111;
		13'b0011000111011: color_data = 12'b010010101111;
		13'b0011000111111: color_data = 12'b010010101111;
		13'b0011001000011: color_data = 12'b010010101111;

		13'b0011010001100: color_data = 12'b010010101111;
		13'b0011010010000: color_data = 12'b010010101111;
		13'b0011010010010: color_data = 12'b010010101111;
		13'b0011010010011: color_data = 12'b010010101111;
		13'b0011010011000: color_data = 12'b010010101111;
		13'b0011010011101: color_data = 12'b010010101111;
		13'b0011010100011: color_data = 12'b010010101111;
		13'b0011010100111: color_data = 12'b010010101111;
		13'b0011010101001: color_data = 12'b010010101111;
		13'b0011010101011: color_data = 12'b010010101111;
		13'b0011010101101: color_data = 12'b010010101111;
		13'b0011010101111: color_data = 12'b010010101111;
		13'b0011010110000: color_data = 12'b010010101111;
		13'b0011010111011: color_data = 12'b010010101111;
		13'b0011010111111: color_data = 12'b010010101111;
		13'b0011011000011: color_data = 12'b010010101111;

		13'b0011100001100: color_data = 12'b010010101111;
		13'b0011100001110: color_data = 12'b010010101111;
		13'b0011100010000: color_data = 12'b010010101111;
		13'b0011100010010: color_data = 12'b010010101111;
		13'b0011100010011: color_data = 12'b010010101111;
		13'b0011100010100: color_data = 12'b010010101111;
		13'b0011100010101: color_data = 12'b010010101111;
		13'b0011100011000: color_data = 12'b010010101111;
		13'b0011100011101: color_data = 12'b010010101111;
		13'b0011100100011: color_data = 12'b010010101111;
		13'b0011100100111: color_data = 12'b010010101111;
		13'b0011100101001: color_data = 12'b010010101111;
		13'b0011100101101: color_data = 12'b010010101111;
		13'b0011100101111: color_data = 12'b010010101111;
		13'b0011100110000: color_data = 12'b010010101111;
		13'b0011100110001: color_data = 12'b010010101111;
		13'b0011100110010: color_data = 12'b010010101111;
		13'b0011100111011: color_data = 12'b010010101111;
		13'b0011100111111: color_data = 12'b010010101111;
		13'b0011101000011: color_data = 12'b010010101111;

		13'b0011110001100: color_data = 12'b010010101111;
		13'b0011110001101: color_data = 12'b010010101111;
		13'b0011110001110: color_data = 12'b010010101111;
		13'b0011110001111: color_data = 12'b010010101111;
		13'b0011110010000: color_data = 12'b010010101111;
		13'b0011110010010: color_data = 12'b010010101111;
		13'b0011110010011: color_data = 12'b010010101111;
		13'b0011110011000: color_data = 12'b010010101111;
		13'b0011110011101: color_data = 12'b010010101111;
		13'b0011110100011: color_data = 12'b010010101111;
		13'b0011110100111: color_data = 12'b010010101111;
		13'b0011110101001: color_data = 12'b010010101111;
		13'b0011110101101: color_data = 12'b010010101111;
		13'b0011110101111: color_data = 12'b010010101111;
		13'b0011110110000: color_data = 12'b010010101111;
		13'b0011110111011: color_data = 12'b010010101111;
		13'b0011110111111: color_data = 12'b010010101111;
		13'b0011111000011: color_data = 12'b010010101111;

		13'b0100000001100: color_data = 12'b010010101111;
		13'b0100000001101: color_data = 12'b010010101111;
		13'b0100000001111: color_data = 12'b010010101111;
		13'b0100000010000: color_data = 12'b010010101111;
		13'b0100000010010: color_data = 12'b010010101111;
		13'b0100000010011: color_data = 12'b010010101111;
		13'b0100000011000: color_data = 12'b010010101111;
		13'b0100000011101: color_data = 12'b010010101111;
		13'b0100000011110: color_data = 12'b010010101111;
		13'b0100000100011: color_data = 12'b010010101111;
		13'b0100000100111: color_data = 12'b010010101111;
		13'b0100000101001: color_data = 12'b010010101111;
		13'b0100000101101: color_data = 12'b010010101111;
		13'b0100000101111: color_data = 12'b010010101111;
		13'b0100000110000: color_data = 12'b010010101111;
		13'b0100000111011: color_data = 12'b010010101111;
		13'b0100000111111: color_data = 12'b010010101111;
		13'b0100001000011: color_data = 12'b010010101111;

		13'b0100010001100: color_data = 12'b010010101111;
		13'b0100010010000: color_data = 12'b010010101111;
		13'b0100010010010: color_data = 12'b010010101111;
		13'b0100010010011: color_data = 12'b010010101111;
		13'b0100010011000: color_data = 12'b010010101111;
		13'b0100010011110: color_data = 12'b010010101111;
		13'b0100010011111: color_data = 12'b010010101111;
		13'b0100010100100: color_data = 12'b010010101111;
		13'b0100010100110: color_data = 12'b010010101111;
		13'b0100010101001: color_data = 12'b010010101111;
		13'b0100010101101: color_data = 12'b010010101111;
		13'b0100010101111: color_data = 12'b010010101111;
		13'b0100010110000: color_data = 12'b010010101111;
		13'b0100010111011: color_data = 12'b010010101111;
		13'b0100011000000: color_data = 12'b010010101111;
		13'b0100011000010: color_data = 12'b010010101111;

		13'b0100100001100: color_data = 12'b010010101111;
		13'b0100100010000: color_data = 12'b010010101111;
		13'b0100100010011: color_data = 12'b010010101111;
		13'b0100100010100: color_data = 12'b010010101111;
		13'b0100100010101: color_data = 12'b010010101111;
		13'b0100100010110: color_data = 12'b010010101111;
		13'b0100100011000: color_data = 12'b010010101111;
		13'b0100100011001: color_data = 12'b010010101111;
		13'b0100100011010: color_data = 12'b010010101111;
		13'b0100100011011: color_data = 12'b010010101111;
		13'b0100100011111: color_data = 12'b010010101111;
		13'b0100100100000: color_data = 12'b010010101111;
		13'b0100100100001: color_data = 12'b010010101111;
		13'b0100100100100: color_data = 12'b010010101111;
		13'b0100100100101: color_data = 12'b010010101111;
		13'b0100100100110: color_data = 12'b010010101111;
		13'b0100100101001: color_data = 12'b010010101111;
		13'b0100100101101: color_data = 12'b010010101111;
		13'b0100100110000: color_data = 12'b010010101111;
		13'b0100100110001: color_data = 12'b010010101111;
		13'b0100100110010: color_data = 12'b010010101111;
		13'b0100100110011: color_data = 12'b010010101111;
		13'b0100100111011: color_data = 12'b010010101111;
		13'b0100101000000: color_data = 12'b010010101111;
		13'b0100101000001: color_data = 12'b010010101111;
		13'b0100101000010: color_data = 12'b010010101111;







		13'b0110010001110: color_data = 12'b101100110101;
		13'b0110010001111: color_data = 12'b101100110101;
		13'b0110010010000: color_data = 12'b101100110101;
		13'b0110010010001: color_data = 12'b101100110101;
		13'b0110010010011: color_data = 12'b101100110101;
		13'b0110010010111: color_data = 12'b101100110101;
		13'b0110010011010: color_data = 12'b101100110101;
		13'b0110010011011: color_data = 12'b101100110101;
		13'b0110010011100: color_data = 12'b101100110101;
		13'b0110010011111: color_data = 12'b101100110101;
		13'b0110010100011: color_data = 12'b101100110101;
		13'b0110010100110: color_data = 12'b101100110101;
		13'b0110010100111: color_data = 12'b101100110101;
		13'b0110010101000: color_data = 12'b101100110101;
		13'b0110010101001: color_data = 12'b101100110101;
		13'b0110010101110: color_data = 12'b101100110101;
		13'b0110010101111: color_data = 12'b101100110101;
		13'b0110010110000: color_data = 12'b101100110101;
		13'b0110010110011: color_data = 12'b101100110101;
		13'b0110010110100: color_data = 12'b101100110101;
		13'b0110010110101: color_data = 12'b101100110101;
		13'b0110010111000: color_data = 12'b101100110101;
		13'b0110010111100: color_data = 12'b101100110101;
		13'b0110010111111: color_data = 12'b101100110101;
		13'b0110011000000: color_data = 12'b101100110101;
		13'b0110011000001: color_data = 12'b101100110101;
		13'b0110011000010: color_data = 12'b101100110101;

		13'b0110100001101: color_data = 12'b101100110101;
		13'b0110100010011: color_data = 12'b101100110101;
		13'b0110100010100: color_data = 12'b101100110101;
		13'b0110100010111: color_data = 12'b101100110101;
		13'b0110100011001: color_data = 12'b101100110101;
		13'b0110100011010: color_data = 12'b101100110101;
		13'b0110100011100: color_data = 12'b101100110101;
		13'b0110100011101: color_data = 12'b101100110101;
		13'b0110100011111: color_data = 12'b101100110101;
		13'b0110100100011: color_data = 12'b101100110101;
		13'b0110100100101: color_data = 12'b101100110101;
		13'b0110100100110: color_data = 12'b101100110101;
		13'b0110100101101: color_data = 12'b101100110101;
		13'b0110100101110: color_data = 12'b101100110101;
		13'b0110100110010: color_data = 12'b101100110101;
		13'b0110100110011: color_data = 12'b101100110101;
		13'b0110100110101: color_data = 12'b101100110101;
		13'b0110100110110: color_data = 12'b101100110101;
		13'b0110100111000: color_data = 12'b101100110101;
		13'b0110100111001: color_data = 12'b101100110101;
		13'b0110100111011: color_data = 12'b101100110101;
		13'b0110100111100: color_data = 12'b101100110101;
		13'b0110100111110: color_data = 12'b101100110101;
		13'b0110100111111: color_data = 12'b101100110101;

		13'b0110110001101: color_data = 12'b101100110101;
		13'b0110110010011: color_data = 12'b101100110101;
		13'b0110110010100: color_data = 12'b101100110101;
		13'b0110110010111: color_data = 12'b101100110101;
		13'b0110110011001: color_data = 12'b101100110101;
		13'b0110110011010: color_data = 12'b101100110101;
		13'b0110110011100: color_data = 12'b101100110101;
		13'b0110110011101: color_data = 12'b101100110101;
		13'b0110110011111: color_data = 12'b101100110101;
		13'b0110110100010: color_data = 12'b101100110101;
		13'b0110110100101: color_data = 12'b101100110101;
		13'b0110110100110: color_data = 12'b101100110101;
		13'b0110110101101: color_data = 12'b101100110101;
		13'b0110110110010: color_data = 12'b101100110101;
		13'b0110110110011: color_data = 12'b101100110101;
		13'b0110110110101: color_data = 12'b101100110101;
		13'b0110110110110: color_data = 12'b101100110101;
		13'b0110110111000: color_data = 12'b101100110101;
		13'b0110110111001: color_data = 12'b101100110101;
		13'b0110110111011: color_data = 12'b101100110101;
		13'b0110110111100: color_data = 12'b101100110101;
		13'b0110110111110: color_data = 12'b101100110101;
		13'b0110110111111: color_data = 12'b101100110101;

		13'b0111000001101: color_data = 12'b101100110101;
		13'b0111000010011: color_data = 12'b101100110101;
		13'b0111000010100: color_data = 12'b101100110101;
		13'b0111000010101: color_data = 12'b101100110101;
		13'b0111000010111: color_data = 12'b101100110101;
		13'b0111000011001: color_data = 12'b101100110101;
		13'b0111000011101: color_data = 12'b101100110101;
		13'b0111000011111: color_data = 12'b101100110101;
		13'b0111000100001: color_data = 12'b101100110101;
		13'b0111000100101: color_data = 12'b101100110101;
		13'b0111000100110: color_data = 12'b101100110101;
		13'b0111000101101: color_data = 12'b101100110101;
		13'b0111000110010: color_data = 12'b101100110101;
		13'b0111000110110: color_data = 12'b101100110101;
		13'b0111000111000: color_data = 12'b101100110101;
		13'b0111000111010: color_data = 12'b101100110101;
		13'b0111000111100: color_data = 12'b101100110101;
		13'b0111000111110: color_data = 12'b101100110101;
		13'b0111000111111: color_data = 12'b101100110101;

		13'b0111010001110: color_data = 12'b101100110101;
		13'b0111010001111: color_data = 12'b101100110101;
		13'b0111010010000: color_data = 12'b101100110101;
		13'b0111010010011: color_data = 12'b101100110101;
		13'b0111010010100: color_data = 12'b101100110101;
		13'b0111010010101: color_data = 12'b101100110101;
		13'b0111010010111: color_data = 12'b101100110101;
		13'b0111010011001: color_data = 12'b101100110101;
		13'b0111010011101: color_data = 12'b101100110101;
		13'b0111010011111: color_data = 12'b101100110101;
		13'b0111010100000: color_data = 12'b101100110101;
		13'b0111010100101: color_data = 12'b101100110101;
		13'b0111010100110: color_data = 12'b101100110101;
		13'b0111010100111: color_data = 12'b101100110101;
		13'b0111010101000: color_data = 12'b101100110101;
		13'b0111010101101: color_data = 12'b101100110101;
		13'b0111010110010: color_data = 12'b101100110101;
		13'b0111010110110: color_data = 12'b101100110101;
		13'b0111010111000: color_data = 12'b101100110101;
		13'b0111010111100: color_data = 12'b101100110101;
		13'b0111010111110: color_data = 12'b101100110101;
		13'b0111010111111: color_data = 12'b101100110101;
		13'b0111011000000: color_data = 12'b101100110101;
		13'b0111011000001: color_data = 12'b101100110101;

		13'b0111100010001: color_data = 12'b101100110101;
		13'b0111100010011: color_data = 12'b101100110101;
		13'b0111100010101: color_data = 12'b101100110101;
		13'b0111100010110: color_data = 12'b101100110101;
		13'b0111100010111: color_data = 12'b101100110101;
		13'b0111100011001: color_data = 12'b101100110101;
		13'b0111100011010: color_data = 12'b101100110101;
		13'b0111100011011: color_data = 12'b101100110101;
		13'b0111100011100: color_data = 12'b101100110101;
		13'b0111100011101: color_data = 12'b101100110101;
		13'b0111100011111: color_data = 12'b101100110101;
		13'b0111100100001: color_data = 12'b101100110101;
		13'b0111100100101: color_data = 12'b101100110101;
		13'b0111100100110: color_data = 12'b101100110101;
		13'b0111100101101: color_data = 12'b101100110101;
		13'b0111100110000: color_data = 12'b101100110101;
		13'b0111100110010: color_data = 12'b101100110101;
		13'b0111100110011: color_data = 12'b101100110101;
		13'b0111100110100: color_data = 12'b101100110101;
		13'b0111100110101: color_data = 12'b101100110101;
		13'b0111100110110: color_data = 12'b101100110101;
		13'b0111100111000: color_data = 12'b101100110101;
		13'b0111100111100: color_data = 12'b101100110101;
		13'b0111100111110: color_data = 12'b101100110101;
		13'b0111100111111: color_data = 12'b101100110101;

		13'b0111110010001: color_data = 12'b101100110101;
		13'b0111110010011: color_data = 12'b101100110101;
		13'b0111110010110: color_data = 12'b101100110101;
		13'b0111110010111: color_data = 12'b101100110101;
		13'b0111110011001: color_data = 12'b101100110101;
		13'b0111110011101: color_data = 12'b101100110101;
		13'b0111110011111: color_data = 12'b101100110101;
		13'b0111110100010: color_data = 12'b101100110101;
		13'b0111110100101: color_data = 12'b101100110101;
		13'b0111110100110: color_data = 12'b101100110101;
		13'b0111110101101: color_data = 12'b101100110101;
		13'b0111110110000: color_data = 12'b101100110101;
		13'b0111110110010: color_data = 12'b101100110101;
		13'b0111110110110: color_data = 12'b101100110101;
		13'b0111110111000: color_data = 12'b101100110101;
		13'b0111110111100: color_data = 12'b101100110101;
		13'b0111110111110: color_data = 12'b101100110101;
		13'b0111110111111: color_data = 12'b101100110101;

		13'b1000000010001: color_data = 12'b101100110101;
		13'b1000000010011: color_data = 12'b101100110101;
		13'b1000000010110: color_data = 12'b101100110101;
		13'b1000000010111: color_data = 12'b101100110101;
		13'b1000000011001: color_data = 12'b101100110101;
		13'b1000000011101: color_data = 12'b101100110101;
		13'b1000000011111: color_data = 12'b101100110101;
		13'b1000000100011: color_data = 12'b101100110101;
		13'b1000000100101: color_data = 12'b101100110101;
		13'b1000000100110: color_data = 12'b101100110101;
		13'b1000000101101: color_data = 12'b101100110101;
		13'b1000000101110: color_data = 12'b101100110101;
		13'b1000000110000: color_data = 12'b101100110101;
		13'b1000000110010: color_data = 12'b101100110101;
		13'b1000000110110: color_data = 12'b101100110101;
		13'b1000000111000: color_data = 12'b101100110101;
		13'b1000000111100: color_data = 12'b101100110101;
		13'b1000000111110: color_data = 12'b101100110101;
		13'b1000000111111: color_data = 12'b101100110101;

		13'b1000010001101: color_data = 12'b101100110101;
		13'b1000010001110: color_data = 12'b101100110101;
		13'b1000010001111: color_data = 12'b101100110101;
		13'b1000010010000: color_data = 12'b101100110101;
		13'b1000010010011: color_data = 12'b101100110101;
		13'b1000010010111: color_data = 12'b101100110101;
		13'b1000010011001: color_data = 12'b101100110101;
		13'b1000010011101: color_data = 12'b101100110101;
		13'b1000010011111: color_data = 12'b101100110101;
		13'b1000010100011: color_data = 12'b101100110101;
		13'b1000010100110: color_data = 12'b101100110101;
		13'b1000010100111: color_data = 12'b101100110101;
		13'b1000010101000: color_data = 12'b101100110101;
		13'b1000010101001: color_data = 12'b101100110101;
		13'b1000010101110: color_data = 12'b101100110101;
		13'b1000010101111: color_data = 12'b101100110101;
		13'b1000010110000: color_data = 12'b101100110101;
		13'b1000010110010: color_data = 12'b101100110101;
		13'b1000010110110: color_data = 12'b101100110101;
		13'b1000010111000: color_data = 12'b101100110101;
		13'b1000010111100: color_data = 12'b101100110101;
		13'b1000010111111: color_data = 12'b101100110101;
		13'b1000011000000: color_data = 12'b101100110101;
		13'b1000011000001: color_data = 12'b101100110101;
		13'b1000011000010: color_data = 12'b101100110101;





		13'b1001100010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1001100010100: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1001100010101: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1001100010110: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1001100010111: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1001100011000: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1001100011001: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1001100011010: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1001100011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1001100100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1001100100101: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1001100100110: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1001100100111: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1001100101000: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1001100101001: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1001100101010: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1001100101011: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1001100101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1001100110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1001100110110: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1001100110111: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1001100111000: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1001100111001: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1001100111010: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1001100111011: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1001100111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h

		13'b1001110010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1001110011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1001110100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1001110101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1001110110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1001110111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h

		13'b1010000010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1010000010110: color_data = 12'b001110100111;
		13'b1010000010111: color_data = 12'b001110100111;
		13'b1010000011000: color_data = 12'b001110100111;
		13'b1010000011001: color_data = 12'b001110100111;
		13'b1010000011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1010000100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1010000100110: color_data = 12'b111110100101;
		13'b1010000101010: color_data = 12'b111110100101;
		13'b1010000101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1010000110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1010000110111: color_data = 12'b101100110101;
		13'b1010000111010: color_data = 12'b101100110101;
		13'b1010000111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h

		13'b1010010010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1010010010101: color_data = 12'b001110100111;
		13'b1010010010110: color_data = 12'b001110100111;
		13'b1010010011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1010010100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1010010100110: color_data = 12'b111110100101;
		13'b1010010100111: color_data = 12'b111110100101;
		13'b1010010101001: color_data = 12'b111110100101;
		13'b1010010101010: color_data = 12'b111110100101;
		13'b1010010101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1010010110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1010010110111: color_data = 12'b101100110101;
		13'b1010010111010: color_data = 12'b101100110101;
		13'b1010010111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h

		13'b1010100010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1010100010101: color_data = 12'b001110100111;
		13'b1010100010110: color_data = 12'b001110100111;
		13'b1010100011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1010100100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1010100100110: color_data = 12'b111110100101;
		13'b1010100100111: color_data = 12'b111110100101;
		13'b1010100101001: color_data = 12'b111110100101;
		13'b1010100101010: color_data = 12'b111110100101; 
		13'b1010100101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1010100110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1010100110111: color_data = 12'b101100110101;
		13'b1010100111010: color_data = 12'b101100110101;
		13'b1010100111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h

		13'b1010110010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1010110010101: color_data = 12'b001110100111;
		13'b1010110010110: color_data = 12'b001110100111;
		13'b1010110011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1010110100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1010110100110: color_data = 12'b111110100101;
		13'b1010110101000: color_data = 12'b111110100101;
		13'b1010110101010: color_data = 12'b111110100101;
		13'b1010110101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1010110110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1010110110111: color_data = 12'b101100110101;
		13'b1010110111010: color_data = 12'b101100110101;
		13'b1010110111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h

		13'b1011000010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1011000010101: color_data = 12'b001110100111;
		13'b1011000010110: color_data = 12'b001110100111;
		13'b1011000010111: color_data = 12'b001110100111;
		13'b1011000011000: color_data = 12'b001110100111;
		13'b1011000011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1011000100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1011000100110: color_data = 12'b111110100101;
		13'b1011000101010: color_data = 12'b111110100101;
		13'b1011000101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1011000110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1011000110111: color_data = 12'b101100110101;
		13'b1011000111000: color_data = 12'b101100110101;
		13'b1011000111001: color_data = 12'b101100110101;
		13'b1011000111010: color_data = 12'b101100110101;
		13'b1011000111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h

		13'b1011010010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1011010010101: color_data = 12'b001110100111;
		13'b1011010010110: color_data = 12'b001110100111;
		13'b1011010011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1011010100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1011010100110: color_data = 12'b111110100101;
		13'b1011010101010: color_data = 12'b111110100101;
		13'b1011010101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1011010110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1011010110111: color_data = 12'b101100110101;
		13'b1011010111010: color_data = 12'b101100110101;
		13'b1011010111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h

		13'b1011100010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e 
		13'b1011100010101: color_data = 12'b001110100111;
		13'b1011100010110: color_data = 12'b001110100111;
		13'b1011100011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1011100100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1011100100110: color_data = 12'b111110100101;
		13'b1011100101010: color_data = 12'b111110100101;
		13'b1011100101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1011100110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1011100110111: color_data = 12'b101100110101;
		13'b1011100111010: color_data = 12'b101100110101;
		13'b1011100111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h

		13'b1011110010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1011110010101: color_data = 12'b001110100111;
		13'b1011110010110: color_data = 12'b001110100111;
		13'b1011110011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1011110100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1011110100110: color_data = 12'b111110100101;
		13'b1011110101010: color_data = 12'b111110100101;
		13'b1011110101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1011110110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1011110110111: color_data = 12'b101100110101;
		13'b1011110111010: color_data = 12'b101100110101;
		13'b1011110111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h

		13'b1100000010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1100000010110: color_data = 12'b001110100111;
		13'b1100000010111: color_data = 12'b001110100111;
		13'b1100000011000: color_data = 12'b001110100111;
		13'b1100000011001: color_data = 12'b001110100111;
		13'b1100000011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1100000100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1100000100110: color_data = 12'b111110100101;
		13'b1100000101010: color_data = 12'b111110100101;
		13'b1100000101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1100000110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1100000110111: color_data = 12'b101100110101;
		13'b1100000111010: color_data = 12'b101100110101;
		13'b1100000111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h

		13'b1100010010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1100010011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1100010100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1100010101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1100010110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1100010111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h

		13'b1100100010011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1100100010100: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1100100010101: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1100100010110: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1100100010111: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1100100011000: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1100100011001: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1100100011010: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		13'b1100100011011: color_data = (mode==2'b00)?12'b111111111111:12'b0; // e
		
		13'b1100100100100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1100100100101: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1100100100110: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1100100100111: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1100100101000: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1100100101001: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1100100101010: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1100100101011: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		13'b1100100101100: color_data = (mode==2'b01)?12'b111111111111:12'b0; // m
		
		13'b1100100110101: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1100100110110: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1100100110111: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1100100111000: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1100100111001: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1100100111010: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1100100111011: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h
		13'b1100100111100: color_data = (mode==2'b10)?12'b111111111111:12'b0; // h 
		default: color_data = 12'b000000000000;
	endcase
endmodule
