`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/28/2025 12:49:25 PM
// Design Name: 
// Module Name: gameOver
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module gameOver(
		input wire clk,
		input wire [4:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})








		11'b01000001100: color_data = 12'b111000010010;
		11'b01000001101: color_data = 12'b111000010010;
		11'b01000001110: color_data = 12'b111000010010;
		11'b01000010001: color_data = 12'b111000010010;
		11'b01000010010: color_data = 12'b111000010010;
		11'b01000010101: color_data = 12'b111000010010;
		11'b01000011000: color_data = 12'b111000010010;
		11'b01000011011: color_data = 12'b111000010010;
		11'b01000011100: color_data = 12'b111000010010;
		11'b01000011101: color_data = 12'b111000010010;

		11'b01001001011: color_data = 12'b111000010010;
		11'b01001010000: color_data = 12'b111000010010;
		11'b01001010011: color_data = 12'b111000010010;
		11'b01001010101: color_data = 12'b111000010010;
		11'b01001010110: color_data = 12'b111000010010;
		11'b01001010111: color_data = 12'b111000010010;
		11'b01001011000: color_data = 12'b111000010010;
		11'b01001011010: color_data = 12'b111000010010;

		11'b01010001011: color_data = 12'b111000010010;
		11'b01010010000: color_data = 12'b111000010010;
		11'b01010010011: color_data = 12'b111000010010;
		11'b01010010101: color_data = 12'b111000010010;
		11'b01010011000: color_data = 12'b111000010010;
		11'b01010011010: color_data = 12'b111000010010;

		11'b01011001011: color_data = 12'b111000010010;
		11'b01011001101: color_data = 12'b111000010010;
		11'b01011001110: color_data = 12'b111000010010;
		11'b01011010000: color_data = 12'b111000010010;
		11'b01011010001: color_data = 12'b111000010010;
		11'b01011010010: color_data = 12'b111000010010;
		11'b01011010011: color_data = 12'b111000010010;
		11'b01011010101: color_data = 12'b111000010010;
		11'b01011011000: color_data = 12'b111000010010;
		11'b01011011010: color_data = 12'b111000010010;
		11'b01011011011: color_data = 12'b111000010010;
		11'b01011011100: color_data = 12'b111000010010;

		11'b01100001011: color_data = 12'b111000010010;
		11'b01100001110: color_data = 12'b111000010010;
		11'b01100010000: color_data = 12'b111000010010;
		11'b01100010011: color_data = 12'b111000010010;
		11'b01100010101: color_data = 12'b111000010010;
		11'b01100011000: color_data = 12'b111000010010;
		11'b01100011010: color_data = 12'b111000010010;

		11'b01101001100: color_data = 12'b111000010010;
		11'b01101001101: color_data = 12'b111000010010;
		11'b01101010000: color_data = 12'b111000010010;
		11'b01101010011: color_data = 12'b111000010010;
		11'b01101010101: color_data = 12'b111000010010;
		11'b01101011000: color_data = 12'b111000010010;
		11'b01101011011: color_data = 12'b111000010010;
		11'b01101011100: color_data = 12'b111000010010;
		11'b01101011101: color_data = 12'b111000010010;



		11'b10000001100: color_data = 12'b111000010010;
		11'b10000001101: color_data = 12'b111000010010;
		11'b10000010000: color_data = 12'b111000010010;
		11'b10000010011: color_data = 12'b111000010010;
		11'b10000010110: color_data = 12'b111000010010;
		11'b10000010111: color_data = 12'b111000010010;
		11'b10000011000: color_data = 12'b111000010010;
		11'b10000011011: color_data = 12'b111000010010;
		11'b10000011100: color_data = 12'b111000010010;

		11'b10001001011: color_data = 12'b111000010010;
		11'b10001001110: color_data = 12'b111000010010;
		11'b10001010000: color_data = 12'b111000010010;
		11'b10001010011: color_data = 12'b111000010010;
		11'b10001010101: color_data = 12'b111000010010;
		11'b10001011010: color_data = 12'b111000010010;
		11'b10001011101: color_data = 12'b111000010010;

		11'b10010001011: color_data = 12'b111000010010;
		11'b10010001110: color_data = 12'b111000010010;
		11'b10010010000: color_data = 12'b111000010010;
		11'b10010010011: color_data = 12'b111000010010;
		11'b10010010101: color_data = 12'b111000010010;
		11'b10010011010: color_data = 12'b111000010010;
		11'b10010011101: color_data = 12'b111000010010;

		11'b10011001011: color_data = 12'b111000010010;
		11'b10011001110: color_data = 12'b111000010010;
		11'b10011010000: color_data = 12'b111000010010;
		11'b10011010011: color_data = 12'b111000010010;
		11'b10011010101: color_data = 12'b111000010010;
		11'b10011010110: color_data = 12'b111000010010;
		11'b10011010111: color_data = 12'b111000010010;
		11'b10011011010: color_data = 12'b111000010010;
		11'b10011011011: color_data = 12'b111000010010;
		11'b10011011100: color_data = 12'b111000010010;

		11'b10100001011: color_data = 12'b111000010010;
		11'b10100001110: color_data = 12'b111000010010;
		11'b10100010000: color_data = 12'b111000010010;
		11'b10100010011: color_data = 12'b111000010010;
		11'b10100010101: color_data = 12'b111000010010;
		11'b10100011010: color_data = 12'b111000010010;
		11'b10100011100: color_data = 12'b111000010010;

		11'b10101001100: color_data = 12'b111000010010;
		11'b10101001101: color_data = 12'b111000010010;
		11'b10101010001: color_data = 12'b111000010010;
		11'b10101010010: color_data = 12'b111000010010;
		11'b10101010110: color_data = 12'b111000010010;
		11'b10101010111: color_data = 12'b111000010010;
		11'b10101011000: color_data = 12'b111000010010;
		11'b10101011010: color_data = 12'b111000010010;
		11'b10101011100: color_data = 12'b111000010010;
		11'b10101011101: color_data = 12'b111000010010;




		default: color_data = 12'b000000000000;
	endcase
endmodule
